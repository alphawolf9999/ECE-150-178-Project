// unsaved_Nios2_A.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module unsaved_Nios2_A (
		output wire [6:0]  HEX_0_external_connection_export,               //              HEX_0_external_connection.export
		output wire [6:0]  HEX_1_external_connection_export,               //              HEX_1_external_connection.export
		output wire [6:0]  HEX_2_external_connection_export,               //              HEX_2_external_connection.export
		output wire [6:0]  HEX_3_external_connection_export,               //              HEX_3_external_connection.export
		output wire [6:0]  HEX_4_external_connection_export,               //              HEX_4_external_connection.export
		output wire [6:0]  HEX_5_external_connection_export,               //              HEX_5_external_connection.export
		output wire [6:0]  HEX_6_external_connection_export,               //              HEX_6_external_connection.export
		output wire [6:0]  HEX_7_external_connection_export,               //              HEX_7_external_connection.export
		output wire [7:0]  LEDG_external_connection_export,                //               LEDG_external_connection.export
		output wire [17:0] LEDR_external_connection_export,                //               LEDR_external_connection.export
		output wire [31:0] avalon_aes_interface_0_export_data_export_data, //     avalon_aes_interface_0_export_data.export_data
		input  wire        clk_0_clk_in_clk,                               //                           clk_0_clk_in.clk
		input  wire        clk_0_clk_in_reset_reset_n,                     //                     clk_0_clk_in_reset.reset_n
		input  wire [3:0]  key_external_connection_export,                 //                key_external_connection.export
		output wire        nios2_gen2_0_custom_instruction_master_readra,  // nios2_gen2_0_custom_instruction_master.readra
		output wire [12:0] sdram_wire_addr,                                //                             sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                                  //                                       .ba
		output wire        sdram_wire_cas_n,                               //                                       .cas_n
		output wire        sdram_wire_cke,                                 //                                       .cke
		output wire        sdram_wire_cs_n,                                //                                       .cs_n
		inout  wire [31:0] sdram_wire_dq,                                  //                                       .dq
		output wire [3:0]  sdram_wire_dqm,                                 //                                       .dqm
		output wire        sdram_wire_ras_n,                               //                                       .ras_n
		output wire        sdram_wire_we_n,                                //                                       .we_n
		input  wire [17:0] switches_external_connection_export             //           switches_external_connection.export
	);

	wire  [31:0] nios2_gen2_0_data_master_readdata;                             // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                          // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                          // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [28:0] nios2_gen2_0_data_master_address;                              // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                           // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                                 // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_readdatavalid;                        // mm_interconnect_0:nios2_gen2_0_data_master_readdatavalid -> nios2_gen2_0:d_readdatavalid
	wire         nios2_gen2_0_data_master_write;                                // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                            // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                      // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                   // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [28:0] nios2_gen2_0_instruction_master_address;                       // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                          // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         nios2_gen2_0_instruction_master_readdatavalid;                 // mm_interconnect_0:nios2_gen2_0_instruction_master_readdatavalid -> nios2_gen2_0:i_readdatavalid
	wire         mm_interconnect_0_avalon_aes_interface_0_aes_slave_chipselect; // mm_interconnect_0:avalon_aes_interface_0_AES_Slave_chipselect -> avalon_aes_interface_0:AVL_CS
	wire  [31:0] mm_interconnect_0_avalon_aes_interface_0_aes_slave_readdata;   // avalon_aes_interface_0:AVL_READDATA -> mm_interconnect_0:avalon_aes_interface_0_AES_Slave_readdata
	wire   [3:0] mm_interconnect_0_avalon_aes_interface_0_aes_slave_address;    // mm_interconnect_0:avalon_aes_interface_0_AES_Slave_address -> avalon_aes_interface_0:AVL_ADDR
	wire         mm_interconnect_0_avalon_aes_interface_0_aes_slave_read;       // mm_interconnect_0:avalon_aes_interface_0_AES_Slave_read -> avalon_aes_interface_0:AVL_READ
	wire   [3:0] mm_interconnect_0_avalon_aes_interface_0_aes_slave_byteenable; // mm_interconnect_0:avalon_aes_interface_0_AES_Slave_byteenable -> avalon_aes_interface_0:AVL_BYTE_EN
	wire         mm_interconnect_0_avalon_aes_interface_0_aes_slave_write;      // mm_interconnect_0:avalon_aes_interface_0_AES_Slave_write -> avalon_aes_interface_0:AVL_WRITE
	wire  [31:0] mm_interconnect_0_avalon_aes_interface_0_aes_slave_writedata;  // mm_interconnect_0:avalon_aes_interface_0_AES_Slave_writedata -> avalon_aes_interface_0:AVL_WRITEDATA
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;    // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;      // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;   // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;          // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;         // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;         // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;          // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;       // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;    // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;    // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;           // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;     // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;          // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;      // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_timer_0_s1_chipselect;                       // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                         // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                          // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                            // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                        // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         mm_interconnect_0_ledr_s1_chipselect;                          // mm_interconnect_0:LEDR_s1_chipselect -> LEDR:chipselect
	wire  [31:0] mm_interconnect_0_ledr_s1_readdata;                            // LEDR:readdata -> mm_interconnect_0:LEDR_s1_readdata
	wire   [1:0] mm_interconnect_0_ledr_s1_address;                             // mm_interconnect_0:LEDR_s1_address -> LEDR:address
	wire         mm_interconnect_0_ledr_s1_write;                               // mm_interconnect_0:LEDR_s1_write -> LEDR:write_n
	wire  [31:0] mm_interconnect_0_ledr_s1_writedata;                           // mm_interconnect_0:LEDR_s1_writedata -> LEDR:writedata
	wire         mm_interconnect_0_ledg_s1_chipselect;                          // mm_interconnect_0:LEDG_s1_chipselect -> LEDG:chipselect
	wire  [31:0] mm_interconnect_0_ledg_s1_readdata;                            // LEDG:readdata -> mm_interconnect_0:LEDG_s1_readdata
	wire   [1:0] mm_interconnect_0_ledg_s1_address;                             // mm_interconnect_0:LEDG_s1_address -> LEDG:address
	wire         mm_interconnect_0_ledg_s1_write;                               // mm_interconnect_0:LEDG_s1_write -> LEDG:write_n
	wire  [31:0] mm_interconnect_0_ledg_s1_writedata;                           // mm_interconnect_0:LEDG_s1_writedata -> LEDG:writedata
	wire         mm_interconnect_0_hex_0_s1_chipselect;                         // mm_interconnect_0:HEX_0_s1_chipselect -> HEX_0:chipselect
	wire  [31:0] mm_interconnect_0_hex_0_s1_readdata;                           // HEX_0:readdata -> mm_interconnect_0:HEX_0_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_0_s1_address;                            // mm_interconnect_0:HEX_0_s1_address -> HEX_0:address
	wire         mm_interconnect_0_hex_0_s1_write;                              // mm_interconnect_0:HEX_0_s1_write -> HEX_0:write_n
	wire  [31:0] mm_interconnect_0_hex_0_s1_writedata;                          // mm_interconnect_0:HEX_0_s1_writedata -> HEX_0:writedata
	wire         mm_interconnect_0_hex_1_s1_chipselect;                         // mm_interconnect_0:HEX_1_s1_chipselect -> HEX_1:chipselect
	wire  [31:0] mm_interconnect_0_hex_1_s1_readdata;                           // HEX_1:readdata -> mm_interconnect_0:HEX_1_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_1_s1_address;                            // mm_interconnect_0:HEX_1_s1_address -> HEX_1:address
	wire         mm_interconnect_0_hex_1_s1_write;                              // mm_interconnect_0:HEX_1_s1_write -> HEX_1:write_n
	wire  [31:0] mm_interconnect_0_hex_1_s1_writedata;                          // mm_interconnect_0:HEX_1_s1_writedata -> HEX_1:writedata
	wire         mm_interconnect_0_hex_2_s1_chipselect;                         // mm_interconnect_0:HEX_2_s1_chipselect -> HEX_2:chipselect
	wire  [31:0] mm_interconnect_0_hex_2_s1_readdata;                           // HEX_2:readdata -> mm_interconnect_0:HEX_2_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_2_s1_address;                            // mm_interconnect_0:HEX_2_s1_address -> HEX_2:address
	wire         mm_interconnect_0_hex_2_s1_write;                              // mm_interconnect_0:HEX_2_s1_write -> HEX_2:write_n
	wire  [31:0] mm_interconnect_0_hex_2_s1_writedata;                          // mm_interconnect_0:HEX_2_s1_writedata -> HEX_2:writedata
	wire         mm_interconnect_0_hex_3_s1_chipselect;                         // mm_interconnect_0:HEX_3_s1_chipselect -> HEX_3:chipselect
	wire  [31:0] mm_interconnect_0_hex_3_s1_readdata;                           // HEX_3:readdata -> mm_interconnect_0:HEX_3_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_3_s1_address;                            // mm_interconnect_0:HEX_3_s1_address -> HEX_3:address
	wire         mm_interconnect_0_hex_3_s1_write;                              // mm_interconnect_0:HEX_3_s1_write -> HEX_3:write_n
	wire  [31:0] mm_interconnect_0_hex_3_s1_writedata;                          // mm_interconnect_0:HEX_3_s1_writedata -> HEX_3:writedata
	wire         mm_interconnect_0_hex_4_s1_chipselect;                         // mm_interconnect_0:HEX_4_s1_chipselect -> HEX_4:chipselect
	wire  [31:0] mm_interconnect_0_hex_4_s1_readdata;                           // HEX_4:readdata -> mm_interconnect_0:HEX_4_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_4_s1_address;                            // mm_interconnect_0:HEX_4_s1_address -> HEX_4:address
	wire         mm_interconnect_0_hex_4_s1_write;                              // mm_interconnect_0:HEX_4_s1_write -> HEX_4:write_n
	wire  [31:0] mm_interconnect_0_hex_4_s1_writedata;                          // mm_interconnect_0:HEX_4_s1_writedata -> HEX_4:writedata
	wire         mm_interconnect_0_hex_5_s1_chipselect;                         // mm_interconnect_0:HEX_5_s1_chipselect -> HEX_5:chipselect
	wire  [31:0] mm_interconnect_0_hex_5_s1_readdata;                           // HEX_5:readdata -> mm_interconnect_0:HEX_5_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_5_s1_address;                            // mm_interconnect_0:HEX_5_s1_address -> HEX_5:address
	wire         mm_interconnect_0_hex_5_s1_write;                              // mm_interconnect_0:HEX_5_s1_write -> HEX_5:write_n
	wire  [31:0] mm_interconnect_0_hex_5_s1_writedata;                          // mm_interconnect_0:HEX_5_s1_writedata -> HEX_5:writedata
	wire         mm_interconnect_0_hex_6_s1_chipselect;                         // mm_interconnect_0:HEX_6_s1_chipselect -> HEX_6:chipselect
	wire  [31:0] mm_interconnect_0_hex_6_s1_readdata;                           // HEX_6:readdata -> mm_interconnect_0:HEX_6_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_6_s1_address;                            // mm_interconnect_0:HEX_6_s1_address -> HEX_6:address
	wire         mm_interconnect_0_hex_6_s1_write;                              // mm_interconnect_0:HEX_6_s1_write -> HEX_6:write_n
	wire  [31:0] mm_interconnect_0_hex_6_s1_writedata;                          // mm_interconnect_0:HEX_6_s1_writedata -> HEX_6:writedata
	wire         mm_interconnect_0_hex_7_s1_chipselect;                         // mm_interconnect_0:HEX_7_s1_chipselect -> HEX_7:chipselect
	wire  [31:0] mm_interconnect_0_hex_7_s1_readdata;                           // HEX_7:readdata -> mm_interconnect_0:HEX_7_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_7_s1_address;                            // mm_interconnect_0:HEX_7_s1_address -> HEX_7:address
	wire         mm_interconnect_0_hex_7_s1_write;                              // mm_interconnect_0:HEX_7_s1_write -> HEX_7:write_n
	wire  [31:0] mm_interconnect_0_hex_7_s1_writedata;                          // mm_interconnect_0:HEX_7_s1_writedata -> HEX_7:writedata
	wire  [31:0] mm_interconnect_0_switches_s1_readdata;                        // switches:readdata -> mm_interconnect_0:switches_s1_readdata
	wire   [1:0] mm_interconnect_0_switches_s1_address;                         // mm_interconnect_0:switches_s1_address -> switches:address
	wire         mm_interconnect_0_highres_s1_chipselect;                       // mm_interconnect_0:highres_s1_chipselect -> highres:chipselect
	wire  [15:0] mm_interconnect_0_highres_s1_readdata;                         // highres:readdata -> mm_interconnect_0:highres_s1_readdata
	wire   [2:0] mm_interconnect_0_highres_s1_address;                          // mm_interconnect_0:highres_s1_address -> highres:address
	wire         mm_interconnect_0_highres_s1_write;                            // mm_interconnect_0:highres_s1_write -> highres:write_n
	wire  [15:0] mm_interconnect_0_highres_s1_writedata;                        // mm_interconnect_0:highres_s1_writedata -> highres:writedata
	wire         mm_interconnect_0_key_s1_chipselect;                           // mm_interconnect_0:key_s1_chipselect -> key:chipselect
	wire  [31:0] mm_interconnect_0_key_s1_readdata;                             // key:readdata -> mm_interconnect_0:key_s1_readdata
	wire   [1:0] mm_interconnect_0_key_s1_address;                              // mm_interconnect_0:key_s1_address -> key:address
	wire         mm_interconnect_0_key_s1_write;                                // mm_interconnect_0:key_s1_write -> key:write_n
	wire  [31:0] mm_interconnect_0_key_s1_writedata;                            // mm_interconnect_0:key_s1_writedata -> key:writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                         // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [31:0] mm_interconnect_0_sdram_s1_readdata;                           // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                        // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                            // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                               // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_s1_byteenable;                         // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                      // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                              // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_s1_writedata;                          // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         irq_mapper_receiver0_irq;                                      // timer_0:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                      // jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                      // key:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                      // highres:irq -> irq_mapper:receiver3_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                          // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                                // rst_controller:reset_out -> [HEX_0:reset_n, HEX_1:reset_n, HEX_2:reset_n, HEX_3:reset_n, HEX_4:reset_n, HEX_5:reset_n, HEX_6:reset_n, HEX_7:reset_n, LEDG:reset_n, LEDR:reset_n, avalon_aes_interface_0:RESET, highres:reset_n, irq_mapper:reset, key:reset_n, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, rst_translator:in_reset, sdram:reset_n, switches:reset_n, sysid_qsys_0:reset_n, timer_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                            // rst_controller:reset_req -> [nios2_gen2_0:reset_req, rst_translator:reset_req_in]
	wire         nios2_gen2_0_debug_reset_request_reset;                        // nios2_gen2_0:debug_reset_request -> [rst_controller:reset_in0, rst_controller_001:reset_in1]
	wire         rst_controller_001_reset_out_reset;                            // rst_controller_001:reset_out -> [jtag_uart_0:rst_n, mm_interconnect_0:jtag_uart_0_reset_reset_bridge_in_reset_reset]

	unsaved_Nios2_A_HEX_0 hex_0 (
		.clk        (clk_0_clk_in_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_0_s1_readdata),   //                    .readdata
		.out_port   (HEX_0_external_connection_export)       // external_connection.export
	);

	unsaved_Nios2_A_HEX_0 hex_1 (
		.clk        (clk_0_clk_in_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_1_s1_readdata),   //                    .readdata
		.out_port   (HEX_1_external_connection_export)       // external_connection.export
	);

	unsaved_Nios2_A_HEX_0 hex_2 (
		.clk        (clk_0_clk_in_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_2_s1_readdata),   //                    .readdata
		.out_port   (HEX_2_external_connection_export)       // external_connection.export
	);

	unsaved_Nios2_A_HEX_0 hex_3 (
		.clk        (clk_0_clk_in_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_3_s1_readdata),   //                    .readdata
		.out_port   (HEX_3_external_connection_export)       // external_connection.export
	);

	unsaved_Nios2_A_HEX_0 hex_4 (
		.clk        (clk_0_clk_in_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_4_s1_readdata),   //                    .readdata
		.out_port   (HEX_4_external_connection_export)       // external_connection.export
	);

	unsaved_Nios2_A_HEX_0 hex_5 (
		.clk        (clk_0_clk_in_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_5_s1_readdata),   //                    .readdata
		.out_port   (HEX_5_external_connection_export)       // external_connection.export
	);

	unsaved_Nios2_A_HEX_0 hex_6 (
		.clk        (clk_0_clk_in_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_6_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_6_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_6_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_6_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_6_s1_readdata),   //                    .readdata
		.out_port   (HEX_6_external_connection_export)       // external_connection.export
	);

	unsaved_Nios2_A_HEX_0 hex_7 (
		.clk        (clk_0_clk_in_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_7_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_7_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_7_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_7_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_7_s1_readdata),   //                    .readdata
		.out_port   (HEX_7_external_connection_export)       // external_connection.export
	);

	unsaved_Nios2_A_LEDG ledg (
		.clk        (clk_0_clk_in_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_ledg_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ledg_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ledg_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ledg_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ledg_s1_readdata),   //                    .readdata
		.out_port   (LEDG_external_connection_export)       // external_connection.export
	);

	unsaved_Nios2_A_LEDR ledr (
		.clk        (clk_0_clk_in_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_ledr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ledr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ledr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ledr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ledr_s1_readdata),   //                    .readdata
		.out_port   (LEDR_external_connection_export)       // external_connection.export
	);

	avalon_aes_interface avalon_aes_interface_0 (
		.RESET         (rst_controller_reset_out_reset),                                //       RESET.reset
		.AVL_CS        (mm_interconnect_0_avalon_aes_interface_0_aes_slave_chipselect), //   AES_Slave.chipselect
		.AVL_BYTE_EN   (mm_interconnect_0_avalon_aes_interface_0_aes_slave_byteenable), //            .byteenable
		.AVL_ADDR      (mm_interconnect_0_avalon_aes_interface_0_aes_slave_address),    //            .address
		.AVL_READ      (mm_interconnect_0_avalon_aes_interface_0_aes_slave_read),       //            .read
		.AVL_READDATA  (mm_interconnect_0_avalon_aes_interface_0_aes_slave_readdata),   //            .readdata
		.AVL_WRITE     (mm_interconnect_0_avalon_aes_interface_0_aes_slave_write),      //            .write
		.AVL_WRITEDATA (mm_interconnect_0_avalon_aes_interface_0_aes_slave_writedata),  //            .writedata
		.EXPORT_DATA   (avalon_aes_interface_0_export_data_export_data),                // Export_Data.export_data
		.CLK           (clk_0_clk_in_clk)                                               //         CLK.clk
	);

	unsaved_Nios2_A_highres highres (
		.clk        (clk_0_clk_in_clk),                        //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_highres_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_highres_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_highres_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_highres_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_highres_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)                 //   irq.irq
	);

	unsaved_Nios2_A_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_0_clk_in_clk),                                            //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                         //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                     //               irq.irq
	);

	unsaved_Nios2_A_key key (
		.clk        (clk_0_clk_in_clk),                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_key_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_key_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_key_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_key_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_key_s1_readdata),   //                    .readdata
		.in_port    (key_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver2_irq)             //                 irq.irq
	);

	unsaved_Nios2_A_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (clk_0_clk_in_clk),                                           //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_gen2_0_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_gen2_0_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       (nios2_gen2_0_custom_instruction_master_readra)               // custom_instruction_master.readra
	);

	unsaved_Nios2_A_sdram sdram (
		.clk            (clk_0_clk_in_clk),                         //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	unsaved_Nios2_A_switches switches (
		.clk      (clk_0_clk_in_clk),                       //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_switches_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_switches_s1_readdata), //                    .readdata
		.in_port  (switches_external_connection_export)     // external_connection.export
	);

	unsaved_Nios2_A_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clk_0_clk_in_clk),                                      //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	unsaved_Nios2_A_timer_0 timer_0 (
		.clk        (clk_0_clk_in_clk),                        //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)                 //   irq.irq
	);

	unsaved_Nios2_A_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                  (clk_0_clk_in_clk),                                              //                                clk_0_clk.clk
		.jtag_uart_0_reset_reset_bridge_in_reset_reset  (rst_controller_001_reset_out_reset),                            //  jtag_uart_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                // nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address               (nios2_gen2_0_data_master_address),                              //                 nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest           (nios2_gen2_0_data_master_waitrequest),                          //                                         .waitrequest
		.nios2_gen2_0_data_master_byteenable            (nios2_gen2_0_data_master_byteenable),                           //                                         .byteenable
		.nios2_gen2_0_data_master_read                  (nios2_gen2_0_data_master_read),                                 //                                         .read
		.nios2_gen2_0_data_master_readdata              (nios2_gen2_0_data_master_readdata),                             //                                         .readdata
		.nios2_gen2_0_data_master_readdatavalid         (nios2_gen2_0_data_master_readdatavalid),                        //                                         .readdatavalid
		.nios2_gen2_0_data_master_write                 (nios2_gen2_0_data_master_write),                                //                                         .write
		.nios2_gen2_0_data_master_writedata             (nios2_gen2_0_data_master_writedata),                            //                                         .writedata
		.nios2_gen2_0_data_master_debugaccess           (nios2_gen2_0_data_master_debugaccess),                          //                                         .debugaccess
		.nios2_gen2_0_instruction_master_address        (nios2_gen2_0_instruction_master_address),                       //          nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest    (nios2_gen2_0_instruction_master_waitrequest),                   //                                         .waitrequest
		.nios2_gen2_0_instruction_master_read           (nios2_gen2_0_instruction_master_read),                          //                                         .read
		.nios2_gen2_0_instruction_master_readdata       (nios2_gen2_0_instruction_master_readdata),                      //                                         .readdata
		.nios2_gen2_0_instruction_master_readdatavalid  (nios2_gen2_0_instruction_master_readdatavalid),                 //                                         .readdatavalid
		.avalon_aes_interface_0_AES_Slave_address       (mm_interconnect_0_avalon_aes_interface_0_aes_slave_address),    //         avalon_aes_interface_0_AES_Slave.address
		.avalon_aes_interface_0_AES_Slave_write         (mm_interconnect_0_avalon_aes_interface_0_aes_slave_write),      //                                         .write
		.avalon_aes_interface_0_AES_Slave_read          (mm_interconnect_0_avalon_aes_interface_0_aes_slave_read),       //                                         .read
		.avalon_aes_interface_0_AES_Slave_readdata      (mm_interconnect_0_avalon_aes_interface_0_aes_slave_readdata),   //                                         .readdata
		.avalon_aes_interface_0_AES_Slave_writedata     (mm_interconnect_0_avalon_aes_interface_0_aes_slave_writedata),  //                                         .writedata
		.avalon_aes_interface_0_AES_Slave_byteenable    (mm_interconnect_0_avalon_aes_interface_0_aes_slave_byteenable), //                                         .byteenable
		.avalon_aes_interface_0_AES_Slave_chipselect    (mm_interconnect_0_avalon_aes_interface_0_aes_slave_chipselect), //                                         .chipselect
		.HEX_0_s1_address                               (mm_interconnect_0_hex_0_s1_address),                            //                                 HEX_0_s1.address
		.HEX_0_s1_write                                 (mm_interconnect_0_hex_0_s1_write),                              //                                         .write
		.HEX_0_s1_readdata                              (mm_interconnect_0_hex_0_s1_readdata),                           //                                         .readdata
		.HEX_0_s1_writedata                             (mm_interconnect_0_hex_0_s1_writedata),                          //                                         .writedata
		.HEX_0_s1_chipselect                            (mm_interconnect_0_hex_0_s1_chipselect),                         //                                         .chipselect
		.HEX_1_s1_address                               (mm_interconnect_0_hex_1_s1_address),                            //                                 HEX_1_s1.address
		.HEX_1_s1_write                                 (mm_interconnect_0_hex_1_s1_write),                              //                                         .write
		.HEX_1_s1_readdata                              (mm_interconnect_0_hex_1_s1_readdata),                           //                                         .readdata
		.HEX_1_s1_writedata                             (mm_interconnect_0_hex_1_s1_writedata),                          //                                         .writedata
		.HEX_1_s1_chipselect                            (mm_interconnect_0_hex_1_s1_chipselect),                         //                                         .chipselect
		.HEX_2_s1_address                               (mm_interconnect_0_hex_2_s1_address),                            //                                 HEX_2_s1.address
		.HEX_2_s1_write                                 (mm_interconnect_0_hex_2_s1_write),                              //                                         .write
		.HEX_2_s1_readdata                              (mm_interconnect_0_hex_2_s1_readdata),                           //                                         .readdata
		.HEX_2_s1_writedata                             (mm_interconnect_0_hex_2_s1_writedata),                          //                                         .writedata
		.HEX_2_s1_chipselect                            (mm_interconnect_0_hex_2_s1_chipselect),                         //                                         .chipselect
		.HEX_3_s1_address                               (mm_interconnect_0_hex_3_s1_address),                            //                                 HEX_3_s1.address
		.HEX_3_s1_write                                 (mm_interconnect_0_hex_3_s1_write),                              //                                         .write
		.HEX_3_s1_readdata                              (mm_interconnect_0_hex_3_s1_readdata),                           //                                         .readdata
		.HEX_3_s1_writedata                             (mm_interconnect_0_hex_3_s1_writedata),                          //                                         .writedata
		.HEX_3_s1_chipselect                            (mm_interconnect_0_hex_3_s1_chipselect),                         //                                         .chipselect
		.HEX_4_s1_address                               (mm_interconnect_0_hex_4_s1_address),                            //                                 HEX_4_s1.address
		.HEX_4_s1_write                                 (mm_interconnect_0_hex_4_s1_write),                              //                                         .write
		.HEX_4_s1_readdata                              (mm_interconnect_0_hex_4_s1_readdata),                           //                                         .readdata
		.HEX_4_s1_writedata                             (mm_interconnect_0_hex_4_s1_writedata),                          //                                         .writedata
		.HEX_4_s1_chipselect                            (mm_interconnect_0_hex_4_s1_chipselect),                         //                                         .chipselect
		.HEX_5_s1_address                               (mm_interconnect_0_hex_5_s1_address),                            //                                 HEX_5_s1.address
		.HEX_5_s1_write                                 (mm_interconnect_0_hex_5_s1_write),                              //                                         .write
		.HEX_5_s1_readdata                              (mm_interconnect_0_hex_5_s1_readdata),                           //                                         .readdata
		.HEX_5_s1_writedata                             (mm_interconnect_0_hex_5_s1_writedata),                          //                                         .writedata
		.HEX_5_s1_chipselect                            (mm_interconnect_0_hex_5_s1_chipselect),                         //                                         .chipselect
		.HEX_6_s1_address                               (mm_interconnect_0_hex_6_s1_address),                            //                                 HEX_6_s1.address
		.HEX_6_s1_write                                 (mm_interconnect_0_hex_6_s1_write),                              //                                         .write
		.HEX_6_s1_readdata                              (mm_interconnect_0_hex_6_s1_readdata),                           //                                         .readdata
		.HEX_6_s1_writedata                             (mm_interconnect_0_hex_6_s1_writedata),                          //                                         .writedata
		.HEX_6_s1_chipselect                            (mm_interconnect_0_hex_6_s1_chipselect),                         //                                         .chipselect
		.HEX_7_s1_address                               (mm_interconnect_0_hex_7_s1_address),                            //                                 HEX_7_s1.address
		.HEX_7_s1_write                                 (mm_interconnect_0_hex_7_s1_write),                              //                                         .write
		.HEX_7_s1_readdata                              (mm_interconnect_0_hex_7_s1_readdata),                           //                                         .readdata
		.HEX_7_s1_writedata                             (mm_interconnect_0_hex_7_s1_writedata),                          //                                         .writedata
		.HEX_7_s1_chipselect                            (mm_interconnect_0_hex_7_s1_chipselect),                         //                                         .chipselect
		.highres_s1_address                             (mm_interconnect_0_highres_s1_address),                          //                               highres_s1.address
		.highres_s1_write                               (mm_interconnect_0_highres_s1_write),                            //                                         .write
		.highres_s1_readdata                            (mm_interconnect_0_highres_s1_readdata),                         //                                         .readdata
		.highres_s1_writedata                           (mm_interconnect_0_highres_s1_writedata),                        //                                         .writedata
		.highres_s1_chipselect                          (mm_interconnect_0_highres_s1_chipselect),                       //                                         .chipselect
		.jtag_uart_0_avalon_jtag_slave_address          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),       //            jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),         //                                         .write
		.jtag_uart_0_avalon_jtag_slave_read             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),          //                                         .read
		.jtag_uart_0_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),      //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),     //                                         .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),   //                                         .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),    //                                         .chipselect
		.key_s1_address                                 (mm_interconnect_0_key_s1_address),                              //                                   key_s1.address
		.key_s1_write                                   (mm_interconnect_0_key_s1_write),                                //                                         .write
		.key_s1_readdata                                (mm_interconnect_0_key_s1_readdata),                             //                                         .readdata
		.key_s1_writedata                               (mm_interconnect_0_key_s1_writedata),                            //                                         .writedata
		.key_s1_chipselect                              (mm_interconnect_0_key_s1_chipselect),                           //                                         .chipselect
		.LEDG_s1_address                                (mm_interconnect_0_ledg_s1_address),                             //                                  LEDG_s1.address
		.LEDG_s1_write                                  (mm_interconnect_0_ledg_s1_write),                               //                                         .write
		.LEDG_s1_readdata                               (mm_interconnect_0_ledg_s1_readdata),                            //                                         .readdata
		.LEDG_s1_writedata                              (mm_interconnect_0_ledg_s1_writedata),                           //                                         .writedata
		.LEDG_s1_chipselect                             (mm_interconnect_0_ledg_s1_chipselect),                          //                                         .chipselect
		.LEDR_s1_address                                (mm_interconnect_0_ledr_s1_address),                             //                                  LEDR_s1.address
		.LEDR_s1_write                                  (mm_interconnect_0_ledr_s1_write),                               //                                         .write
		.LEDR_s1_readdata                               (mm_interconnect_0_ledr_s1_readdata),                            //                                         .readdata
		.LEDR_s1_writedata                              (mm_interconnect_0_ledr_s1_writedata),                           //                                         .writedata
		.LEDR_s1_chipselect                             (mm_interconnect_0_ledr_s1_chipselect),                          //                                         .chipselect
		.nios2_gen2_0_debug_mem_slave_address           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),        //             nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),          //                                         .write
		.nios2_gen2_0_debug_mem_slave_read              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),           //                                         .read
		.nios2_gen2_0_debug_mem_slave_readdata          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),       //                                         .readdata
		.nios2_gen2_0_debug_mem_slave_writedata         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),      //                                         .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),     //                                         .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),    //                                         .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),    //                                         .debugaccess
		.sdram_s1_address                               (mm_interconnect_0_sdram_s1_address),                            //                                 sdram_s1.address
		.sdram_s1_write                                 (mm_interconnect_0_sdram_s1_write),                              //                                         .write
		.sdram_s1_read                                  (mm_interconnect_0_sdram_s1_read),                               //                                         .read
		.sdram_s1_readdata                              (mm_interconnect_0_sdram_s1_readdata),                           //                                         .readdata
		.sdram_s1_writedata                             (mm_interconnect_0_sdram_s1_writedata),                          //                                         .writedata
		.sdram_s1_byteenable                            (mm_interconnect_0_sdram_s1_byteenable),                         //                                         .byteenable
		.sdram_s1_readdatavalid                         (mm_interconnect_0_sdram_s1_readdatavalid),                      //                                         .readdatavalid
		.sdram_s1_waitrequest                           (mm_interconnect_0_sdram_s1_waitrequest),                        //                                         .waitrequest
		.sdram_s1_chipselect                            (mm_interconnect_0_sdram_s1_chipselect),                         //                                         .chipselect
		.switches_s1_address                            (mm_interconnect_0_switches_s1_address),                         //                              switches_s1.address
		.switches_s1_readdata                           (mm_interconnect_0_switches_s1_readdata),                        //                                         .readdata
		.sysid_qsys_0_control_slave_address             (mm_interconnect_0_sysid_qsys_0_control_slave_address),          //               sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata            (mm_interconnect_0_sysid_qsys_0_control_slave_readdata),         //                                         .readdata
		.timer_0_s1_address                             (mm_interconnect_0_timer_0_s1_address),                          //                               timer_0_s1.address
		.timer_0_s1_write                               (mm_interconnect_0_timer_0_s1_write),                            //                                         .write
		.timer_0_s1_readdata                            (mm_interconnect_0_timer_0_s1_readdata),                         //                                         .readdata
		.timer_0_s1_writedata                           (mm_interconnect_0_timer_0_s1_writedata),                        //                                         .writedata
		.timer_0_s1_chipselect                          (mm_interconnect_0_timer_0_s1_chipselect)                        //                                         .chipselect
	);

	unsaved_Nios2_A_irq_mapper irq_mapper (
		.clk           (clk_0_clk_in_clk),               //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.sender_irq    (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (nios2_gen2_0_debug_reset_request_reset), // reset_in0.reset
		.clk            (clk_0_clk_in_clk),                       //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),         // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),     //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~clk_0_clk_in_reset_reset_n),            // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_0_clk_in_clk),                       //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
